library IEEE;
use IEEE.std_logic_1164.all;

entity alu_control is
    port(
        i_ALUOp  : in  std_logic_vector(1 downto 0);  -- From control unit
        i_Funct3 : in  std_logic_vector(2 downto 0);  -- Instruction bits
        i_Funct7 : in  std_logic_vector(6 downto 0);  -- Instruction bits
        o_ALUCtrl: out std_logic_vector(3 downto 0)   -- To ALU
    );
end alu_control;

architecture behavior of alu_control is
begin
    process(i_ALUOp, i_Funct3, i_Funct7)
    begin

        case i_ALUOp is
            --------------------------------------------------------------------
            -- ALUOp = 00 → 기본 ADD (Load, Store, AUIPC)
            --------------------------------------------------------------------
            when "00" =>
                o_ALUCtrl <= "0010";  -- ADD

            --------------------------------------------------------------------
            -- ALUOp = 01 → Branch 연산용 (SUB)
            --------------------------------------------------------------------
            when "01" =>
                o_ALUCtrl <= "0110";  -- SUB

            --------------------------------------------------------------------
            -- ALUOp = 10 → R-type / I-type ALU
            --------------------------------------------------------------------
            when "10" =>
                case i_Funct3 is

                    ----------------------------------------------------------------
                    -- ADD / SUB
                    ----------------------------------------------------------------
                    when "000" =>
                        if i_Funct7 = "0100000" then
                            o_ALUCtrl <= "0110"; -- SUB
                        else
                            o_ALUCtrl <= "0010"; -- ADD / ADDI
                        end if;

                    ----------------------------------------------------------------
                    -- SLL
                    ----------------------------------------------------------------
                    when "001" =>
                        o_ALUCtrl <= "1001"; -- SLL

                    ----------------------------------------------------------------
                    -- SLT
                    ----------------------------------------------------------------
                    when "010" =>
                        o_ALUCtrl <= "0111"; -- SLT
                    
                    ----------------------------------------------------------------
                    -- SLT
                    ----------------------------------------------------------------
                    when "011" =>
                        o_ALUCtrl <= "1100"; -- SLTU/SLTIU

                    ----------------------------------------------------------------
                    -- XOR
                    ----------------------------------------------------------------
                    when "100" =>
                        o_ALUCtrl <= "0100"; -- XOR

                    ----------------------------------------------------------------
                    -- SRL/SRA
                    ----------------------------------------------------------------
                    when "101" =>
                        if i_Funct7 = "0100000" then
                            o_ALUCtrl <= "1010"; -- SRA
                        else
                            o_ALUCtrl <= "1000"; -- SRL
                        end if;

                    ----------------------------------------------------------------
                    -- OR
                    ----------------------------------------------------------------
                    when "110" =>
                        o_ALUCtrl <= "0001"; -- OR

                    ----------------------------------------------------------------
                    -- AND
                    ----------------------------------------------------------------
                    when "111" =>
                        o_ALUCtrl <= "0000"; -- AND

                    when others =>
                        o_ALUCtrl <= "0000";
                end case;
                

            when others =>
                o_ALUCtrl <= "0000";
            

        end case;
    end process;

end behavior;